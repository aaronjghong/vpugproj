logic [TILE_WIDTH-1:0][TILE_HEIGHT-1:0] texture_data_fill [ASCII_LEVELS-1:0] = '{
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 0
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 255, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 1
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 255, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 255, 0, 0, 0},
        '{0, 0, 0, 0, 255, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 2
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 255, 255, 0, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 255, 0, 0, 0, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 0, 255, 255, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 3
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 255, 255, 0, 0, 0, 0},
        '{0, 255, 0, 0, 255, 0, 0, 0},
        '{0, 255, 0, 0, 255, 0, 0, 0},
        '{0, 255, 0, 0, 255, 0, 0, 0},
        '{0, 0, 255, 255, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 4
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 255, 255, 255, 0, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 255, 255, 255, 0, 0, 0},
        '{0, 0, 255, 0, 0, 0, 0, 0},
        '{0, 0, 255, 0, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 5
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 255, 255, 0, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 0, 255, 255, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 6
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 255, 255, 0, 0, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 0, 0, 255, 255, 0, 0},
        '{0, 0, 0, 255, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 255, 0, 0, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 7
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 0, 0, 255, 255, 255, 0, 0},
        '{0, 0, 255, 0, 0, 0, 255, 0},
        '{0, 0, 255, 0, 255, 255, 255, 0},
        '{0, 0, 255, 0, 0, 255, 0, 0},
        '{0, 0, 0, 255, 0, 0, 0, 0},
        '{0, 0, 0, 0, 255, 255, 0, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }, // Character 8
    '{
        '{0, 0, 0, 0, 0, 0, 0, 0},
        '{0, 255, 255, 255, 255, 255, 255, 0},
        '{0, 255, 255, 255, 255, 255, 255, 0},
        '{0, 255, 255, 255, 255, 255, 255, 0},
        '{0, 255, 255, 255, 255, 255, 255, 0},
        '{0, 255, 255, 255, 255, 255, 255, 0},
        '{0, 255, 255, 255, 255, 255, 255, 0},
        '{0, 0, 0, 0, 0, 0, 0, 0}
    }  // Character 9
};
